// Copyright (C) 2020  Intel Corporation. All rights reserved.
// Your use of Intel Corporation's design tools, logic functions 
// and other software and tools, and any partner logic 
// functions, and any output files from any of the foregoing 
// (including device programming or simulation files), and any 
// associated documentation or information are expressly subject 
// to the terms and conditions of the Intel Program License 
// Subscription Agreement, the Intel Quartus Prime License Agreement,
// the Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is for
// the sole purpose of programming logic devices manufactured by
// Intel and sold by Intel or its authorized distributors.  Please
// refer to the applicable agreement for further details, at
// https://fpgasoftware.intel.com/eula.

// Generated by Quartus Prime Version 20.1.0 Build 711 06/05/2020 SJ Lite Edition
// Created on Mon Dec 07 03:59:48 2020

// synthesis message_off 10175

`timescale 1ns/1ns

module SM1 (
    input reset, input clock, input x,
    output y);

    enum int unsigned { state1=0, state2=1, state3=2 } fstate, reg_fstate;

    always_ff @(posedge clock)
    begin
        if (clock) begin
            fstate <= reg_fstate;
        end
    end

    always_comb begin
        if (reset) begin
            reg_fstate <= state1;
            y <= 1'b0;
        end
        else begin
            y <= 1'b0;
            case (fstate)
                state1: begin
                    if ((x == 1'b0))
                        reg_fstate <= state1;
                    else if ((x == 1'b1))
                        reg_fstate <= state2;
                    // Inserting 'else' block to prevent latch inference
                    else
                        reg_fstate <= state1;
                end
                state2: begin
                    if ((x == 1'b1))
                        reg_fstate <= state3;
                    else if ((x == 1'b0))
                        reg_fstate <= state1;
                    // Inserting 'else' block to prevent latch inference
                    else
                        reg_fstate <= state2;
                end
                state3: begin
                    if ((x == 1'b1))
                        reg_fstate <= state3;
                    else if ((x == 1'b0))
                        reg_fstate <= state1;
                    // Inserting 'else' block to prevent latch inference
                    else
                        reg_fstate <= state3;

                    if ((x == 1'b1))
                        y <= 1'b1;
                    // Inserting 'else' block to prevent latch inference
                    else
                        y <= 1'b0;
                end
                default: begin
                    y <= 1'bx;
                    $display ("Reach undefined state");
                end
            endcase
        end
    end
endmodule // SM1
